`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer:    Daniele Ricciardelli
// Design Name: 
// Module Name: incrementer
//////////////////////////////////////////////////////////////////////////////////

module incrementer
(
    input [31:0] pcin,
    output [31:0] pcout     
);
    
    assign pcout = pcin + 32'd4;

endmodule
